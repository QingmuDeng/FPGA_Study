module hello_test ();
initial begin
    $display("hello CompArch");
end
endmodule
